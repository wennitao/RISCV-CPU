`include "cpu_define.v"
// RISCV32I CPU top module
// port modification allowed for debugging purposes
module cpu(
  input  wire                 clk_in,			// system clock signal
  input  wire                 rst_in,			// reset signal
	input  wire					        rdy_in,			// ready signal, pause cpu when low

  input  wire [ 7:0]          mem_din,		// data input bus
  output wire [ 7:0]          mem_dout,		// data output bus
  output wire [31:0]          mem_a,			// address bus (only 17:0 is used)
  output wire                 mem_wr,			// write/read signal (1 for write)
	
	input  wire                 io_buffer_full, // 1 if uart buffer is full
	
	output wire [31:0]			dbgreg_dout		// cpu register output (debugging demo)
);

// implementation goes here

// Specifications:
// - Pause cpu(freeze pc, registers, etc.) when rdy_in is low
// - Memory read result will be returned in the next cycle. Write takes 1 cycle(no need to wait)
// - Memory is of size 128KB, with valid address ranging from 0x0 to 0x20000
// - I/O port is mapped to address higher than 0x30000 (mem_a[17:16]==2'b11)
// - 0x30000 read: read a byte from input
// - 0x30000 write: write a byte to output (write 0x00 is ignored)
// - 0x30004 read: read clocks passed since cpu starts (in dword, 4 bytes)
// - 0x30004 write: indicates program stop (will output '\0' through uart tx)

// MemCtrl <-> InstCache
wire MemCtrl_InstCache_inst_read_valid, MemCtrl_InstCache_inst_valid ;
wire [`AddressBus] MemCtrl_InstCache_inst_addr ;
wire [`InstBus] MemCtrl_InstCache_inst ;

// InstCache <-> IF
wire InstCache_IF_inst_valid, InstCache_IF_inst_read_valid ;
wire [`AddressBus] InstCache_IF_inst_addr ;
wire [`InstBus] InstCache_IF_inst ;

MemCtrl MemCtrl (
  .clk (clk_in), 
  .rst (rst_in), 
  .rdy (rdy_in), 

  .InstCache_inst_read_valid (MemCtrl_InstCache_inst_read_valid), 
  .InstCache_inst_addr (MemCtrl_InstCache_inst_addr), 
  .InstCache_inst_valid (MemCtrl_InstCache_inst_valid), 
  .InstCache_inst (MemCtrl_InstCache_inst), 

  .mem_din (mem_din), 
  .mem_dout (mem_dout), 
  .mem_a (mem_a), 
  .mem_wr (mem_wr)
) ;

InstructionCache InstructionCache (
  .clk (clk_in), 
  .rst (rst_in), 
  .rdy (rdy_in), 

  .IF_inst_read_valid (InstCache_IF_inst_read_valid), 
  .IF_inst_addr (InstCache_IF_inst_addr), 
  .IF_inst_valid (InstCache_IF_inst_valid), 
  .IF_inst (InstCache_IF_inst), 

  .MemCtrl_inst_valid (MemCtrl_InstCache_inst_valid), 
  .MemCtrl_inst (MemCtrl_InstCache_inst), 
  .MemCtrl_inst_read_valid (MemCtrl_InstCache_inst_read_valid), 
  .MemCtrl_inst_addr (MemCtrl_InstCache_inst_addr)
) ;

IF IF (
  .clk (clk_in), 
  .rst (rst_in), 
  .rdy (rdy_in), 

  .InstCache_inst_valid (InstCache_IF_inst_valid), 
  .InstCache_inst (InstCache_IF_inst), 
  .InstCache_inst_read_valid (InstCache_IF_inst_read_valid), 
  .InstCache_inst_addr (InstCache_IF_inst_addr)
) ;

endmodule